//single-precision floating point as defined by IEEE 754
parameter int DATA_WIDTH = 32
parameter int EXPONENT_WIDTH = 8
parameter int MANTISA_WIDTH = 23